`ifndef CONFIG_VH
`define CONFIG_VH

`timescale 1 ns / 1 ps

`define USE_STRUCTURAL_IMPLEMENTATION

// `define CLK_100_MHZ
   `define CLK_50_MHZ
// `define CLK_25_MHZ

`endif
