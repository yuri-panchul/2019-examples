`ifndef GAME_CONFIG_VH
`define GAME_CONFIG_VH

`include "config.vh"

`endif
