module fsm_3_bits_coming_from_left
(
    input        clk,
    input        rst,
    input        new_bit,
    output [1:0] rem
);

    assign rem = 0;

endmodule
